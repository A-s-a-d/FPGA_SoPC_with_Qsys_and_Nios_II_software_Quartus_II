// de1_blinker.v

// Generated using ACDS version 15.0 153

`timescale 1 ps / 1 ps
module de1_blinker (
		output wire [2:0] calibration_external_connection_export, // calibration_external_connection.export
		input  wire [3:0] centaines_external_connection_export,   //   centaines_external_connection.export
		input  wire       clk_clk,                                //                             clk.clk
		input  wire [3:0] dizaines_external_connection_export,    //    dizaines_external_connection.export
		output wire [7:0] led_external_connection_export,         //         led_external_connection.export
		input  wire [3:0] milliers_external_connection_export,    //    milliers_external_connection.export
		output wire [7:0] seven_seg_1_external_connection_export, // seven_seg_1_external_connection.export
		output wire [7:0] seven_seg_2_external_connection_export, // seven_seg_2_external_connection.export
		output wire [7:0] seven_seg_3_external_connection_export, // seven_seg_3_external_connection.export
		output wire [7:0] seven_seg_4_external_connection_export, // seven_seg_4_external_connection.export
		input  wire [3:0] switcher_external_connection_export,    //    switcher_external_connection.export
		input  wire [3:0] unites_external_connection_export       //      unites_external_connection.export
	);

	wire         nios2_proc_jtag_debug_module_reset_reset;                    // nios2_proc:jtag_debug_module_resetrequest -> rst_controller:reset_in0
	wire  [31:0] nios2_proc_data_master_readdata;                             // mm_interconnect_0:nios2_proc_data_master_readdata -> nios2_proc:d_readdata
	wire         nios2_proc_data_master_waitrequest;                          // mm_interconnect_0:nios2_proc_data_master_waitrequest -> nios2_proc:d_waitrequest
	wire         nios2_proc_data_master_debugaccess;                          // nios2_proc:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_proc_data_master_debugaccess
	wire  [19:0] nios2_proc_data_master_address;                              // nios2_proc:d_address -> mm_interconnect_0:nios2_proc_data_master_address
	wire   [3:0] nios2_proc_data_master_byteenable;                           // nios2_proc:d_byteenable -> mm_interconnect_0:nios2_proc_data_master_byteenable
	wire         nios2_proc_data_master_read;                                 // nios2_proc:d_read -> mm_interconnect_0:nios2_proc_data_master_read
	wire         nios2_proc_data_master_write;                                // nios2_proc:d_write -> mm_interconnect_0:nios2_proc_data_master_write
	wire  [31:0] nios2_proc_data_master_writedata;                            // nios2_proc:d_writedata -> mm_interconnect_0:nios2_proc_data_master_writedata
	wire  [31:0] nios2_proc_instruction_master_readdata;                      // mm_interconnect_0:nios2_proc_instruction_master_readdata -> nios2_proc:i_readdata
	wire         nios2_proc_instruction_master_waitrequest;                   // mm_interconnect_0:nios2_proc_instruction_master_waitrequest -> nios2_proc:i_waitrequest
	wire  [19:0] nios2_proc_instruction_master_address;                       // nios2_proc:i_address -> mm_interconnect_0:nios2_proc_instruction_master_address
	wire         nios2_proc_instruction_master_read;                          // nios2_proc:i_read -> mm_interconnect_0:nios2_proc_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_1337_control_slave_readdata;         // sysid_1337:readdata -> mm_interconnect_0:sysid_1337_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_1337_control_slave_address;          // mm_interconnect_0:sysid_1337_control_slave_address -> sysid_1337:address
	wire  [31:0] mm_interconnect_0_nios2_proc_jtag_debug_module_readdata;     // nios2_proc:jtag_debug_module_readdata -> mm_interconnect_0:nios2_proc_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_proc_jtag_debug_module_waitrequest;  // nios2_proc:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_proc_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_proc_jtag_debug_module_debugaccess;  // mm_interconnect_0:nios2_proc_jtag_debug_module_debugaccess -> nios2_proc:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_proc_jtag_debug_module_address;      // mm_interconnect_0:nios2_proc_jtag_debug_module_address -> nios2_proc:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_proc_jtag_debug_module_read;         // mm_interconnect_0:nios2_proc_jtag_debug_module_read -> nios2_proc:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_proc_jtag_debug_module_byteenable;   // mm_interconnect_0:nios2_proc_jtag_debug_module_byteenable -> nios2_proc:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_proc_jtag_debug_module_write;        // mm_interconnect_0:nios2_proc_jtag_debug_module_write -> nios2_proc:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_proc_jtag_debug_module_writedata;    // mm_interconnect_0:nios2_proc_jtag_debug_module_writedata -> nios2_proc:jtag_debug_module_writedata
	wire         mm_interconnect_0_led_s1_chipselect;                         // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                           // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                            // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                              // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                          // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire  [31:0] mm_interconnect_0_switcher_s1_readdata;                      // switcher:readdata -> mm_interconnect_0:switcher_s1_readdata
	wire   [1:0] mm_interconnect_0_switcher_s1_address;                       // mm_interconnect_0:switcher_s1_address -> switcher:address
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;               // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                 // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory_s1_address;                  // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;               // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                    // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                    // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_seven_seg_1_s1_chipselect;                 // mm_interconnect_0:Seven_Seg_1_s1_chipselect -> Seven_Seg_1:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_1_s1_readdata;                   // Seven_Seg_1:readdata -> mm_interconnect_0:Seven_Seg_1_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_1_s1_address;                    // mm_interconnect_0:Seven_Seg_1_s1_address -> Seven_Seg_1:address
	wire         mm_interconnect_0_seven_seg_1_s1_write;                      // mm_interconnect_0:Seven_Seg_1_s1_write -> Seven_Seg_1:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_1_s1_writedata;                  // mm_interconnect_0:Seven_Seg_1_s1_writedata -> Seven_Seg_1:writedata
	wire         mm_interconnect_0_seven_seg_4_s1_chipselect;                 // mm_interconnect_0:Seven_Seg_4_s1_chipselect -> Seven_Seg_4:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_4_s1_readdata;                   // Seven_Seg_4:readdata -> mm_interconnect_0:Seven_Seg_4_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_4_s1_address;                    // mm_interconnect_0:Seven_Seg_4_s1_address -> Seven_Seg_4:address
	wire         mm_interconnect_0_seven_seg_4_s1_write;                      // mm_interconnect_0:Seven_Seg_4_s1_write -> Seven_Seg_4:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_4_s1_writedata;                  // mm_interconnect_0:Seven_Seg_4_s1_writedata -> Seven_Seg_4:writedata
	wire         mm_interconnect_0_seven_seg_3_s1_chipselect;                 // mm_interconnect_0:Seven_Seg_3_s1_chipselect -> Seven_Seg_3:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_3_s1_readdata;                   // Seven_Seg_3:readdata -> mm_interconnect_0:Seven_Seg_3_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_3_s1_address;                    // mm_interconnect_0:Seven_Seg_3_s1_address -> Seven_Seg_3:address
	wire         mm_interconnect_0_seven_seg_3_s1_write;                      // mm_interconnect_0:Seven_Seg_3_s1_write -> Seven_Seg_3:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_3_s1_writedata;                  // mm_interconnect_0:Seven_Seg_3_s1_writedata -> Seven_Seg_3:writedata
	wire         mm_interconnect_0_seven_seg_2_s1_chipselect;                 // mm_interconnect_0:Seven_Seg_2_s1_chipselect -> Seven_Seg_2:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_2_s1_readdata;                   // Seven_Seg_2:readdata -> mm_interconnect_0:Seven_Seg_2_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_2_s1_address;                    // mm_interconnect_0:Seven_Seg_2_s1_address -> Seven_Seg_2:address
	wire         mm_interconnect_0_seven_seg_2_s1_write;                      // mm_interconnect_0:Seven_Seg_2_s1_write -> Seven_Seg_2:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_2_s1_writedata;                  // mm_interconnect_0:Seven_Seg_2_s1_writedata -> Seven_Seg_2:writedata
	wire  [31:0] mm_interconnect_0_unites_s1_readdata;                        // Unites:readdata -> mm_interconnect_0:Unites_s1_readdata
	wire   [1:0] mm_interconnect_0_unites_s1_address;                         // mm_interconnect_0:Unites_s1_address -> Unites:address
	wire  [31:0] mm_interconnect_0_dizaines_s1_readdata;                      // Dizaines:readdata -> mm_interconnect_0:Dizaines_s1_readdata
	wire   [1:0] mm_interconnect_0_dizaines_s1_address;                       // mm_interconnect_0:Dizaines_s1_address -> Dizaines:address
	wire  [31:0] mm_interconnect_0_centaines_s1_readdata;                     // Centaines:readdata -> mm_interconnect_0:Centaines_s1_readdata
	wire   [1:0] mm_interconnect_0_centaines_s1_address;                      // mm_interconnect_0:Centaines_s1_address -> Centaines:address
	wire  [31:0] mm_interconnect_0_milliers_s1_readdata;                      // Milliers:readdata -> mm_interconnect_0:Milliers_s1_readdata
	wire   [1:0] mm_interconnect_0_milliers_s1_address;                       // mm_interconnect_0:Milliers_s1_address -> Milliers:address
	wire         mm_interconnect_0_calibration_s1_chipselect;                 // mm_interconnect_0:Calibration_s1_chipselect -> Calibration:chipselect
	wire  [31:0] mm_interconnect_0_calibration_s1_readdata;                   // Calibration:readdata -> mm_interconnect_0:Calibration_s1_readdata
	wire   [1:0] mm_interconnect_0_calibration_s1_address;                    // mm_interconnect_0:Calibration_s1_address -> Calibration:address
	wire         mm_interconnect_0_calibration_s1_write;                      // mm_interconnect_0:Calibration_s1_write -> Calibration:write_n
	wire  [31:0] mm_interconnect_0_calibration_s1_writedata;                  // mm_interconnect_0:Calibration_s1_writedata -> Calibration:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_proc_d_irq_irq;                                        // irq_mapper:sender_irq -> nios2_proc:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [Calibration:reset_n, Centaines:reset_n, Dizaines:reset_n, Milliers:reset_n, Seven_Seg_1:reset_n, Seven_Seg_2:reset_n, Seven_Seg_3:reset_n, Seven_Seg_4:reset_n, Unites:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, led:reset_n, mm_interconnect_0:nios2_proc_reset_n_reset_bridge_in_reset_reset, nios2_proc:reset_n, onchip_memory:reset, rst_translator:in_reset, switcher:reset_n, sysid_1337:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_proc:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]

	de1_blinker_Calibration calibration (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_calibration_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_calibration_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_calibration_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_calibration_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_calibration_s1_readdata),   //                    .readdata
		.out_port   (calibration_external_connection_export)       // external_connection.export
	);

	de1_blinker_Centaines centaines (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_centaines_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_centaines_s1_readdata), //                    .readdata
		.in_port  (centaines_external_connection_export)     // external_connection.export
	);

	de1_blinker_Centaines dizaines (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_dizaines_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dizaines_s1_readdata), //                    .readdata
		.in_port  (dizaines_external_connection_export)     // external_connection.export
	);

	de1_blinker_Centaines milliers (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_milliers_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_milliers_s1_readdata), //                    .readdata
		.in_port  (milliers_external_connection_export)     // external_connection.export
	);

	de1_blinker_Seven_Seg_1 seven_seg_1 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_1_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_1_external_connection_export)       // external_connection.export
	);

	de1_blinker_Seven_Seg_1 seven_seg_2 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_2_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_2_external_connection_export)       // external_connection.export
	);

	de1_blinker_Seven_Seg_1 seven_seg_3 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_3_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_3_external_connection_export)       // external_connection.export
	);

	de1_blinker_Seven_Seg_1 seven_seg_4 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_4_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_4_external_connection_export)       // external_connection.export
	);

	de1_blinker_Centaines unites (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_unites_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_unites_s1_readdata), //                    .readdata
		.in_port  (unites_external_connection_export)     // external_connection.export
	);

	de1_blinker_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	de1_blinker_Seven_Seg_1 led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	de1_blinker_nios2_proc nios2_proc (
		.clk                                   (clk_clk),                                                    //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                            //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                             (nios2_proc_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_proc_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_proc_data_master_read),                                //                          .read
		.d_readdata                            (nios2_proc_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_proc_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_proc_data_master_write),                               //                          .write
		.d_writedata                           (nios2_proc_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_proc_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_proc_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_proc_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_proc_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_proc_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_proc_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_proc_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_proc_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_proc_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_proc_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_proc_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_proc_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_proc_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_proc_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_proc_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                            // custom_instruction_master.readra
	);

	de1_blinker_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	de1_blinker_Centaines switcher (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switcher_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switcher_s1_readdata), //                    .readdata
		.in_port  (switcher_external_connection_export)     // external_connection.export
	);

	de1_blinker_sysid_1337 sysid_1337 (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_1337_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_1337_control_slave_address)   //              .address
	);

	de1_blinker_mm_interconnect_0 mm_interconnect_0 (
		.clk_main_clk_clk                               (clk_clk),                                                     //                             clk_main_clk.clk
		.nios2_proc_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_proc_reset_n_reset_bridge_in_reset.reset
		.nios2_proc_data_master_address                 (nios2_proc_data_master_address),                              //                   nios2_proc_data_master.address
		.nios2_proc_data_master_waitrequest             (nios2_proc_data_master_waitrequest),                          //                                         .waitrequest
		.nios2_proc_data_master_byteenable              (nios2_proc_data_master_byteenable),                           //                                         .byteenable
		.nios2_proc_data_master_read                    (nios2_proc_data_master_read),                                 //                                         .read
		.nios2_proc_data_master_readdata                (nios2_proc_data_master_readdata),                             //                                         .readdata
		.nios2_proc_data_master_write                   (nios2_proc_data_master_write),                                //                                         .write
		.nios2_proc_data_master_writedata               (nios2_proc_data_master_writedata),                            //                                         .writedata
		.nios2_proc_data_master_debugaccess             (nios2_proc_data_master_debugaccess),                          //                                         .debugaccess
		.nios2_proc_instruction_master_address          (nios2_proc_instruction_master_address),                       //            nios2_proc_instruction_master.address
		.nios2_proc_instruction_master_waitrequest      (nios2_proc_instruction_master_waitrequest),                   //                                         .waitrequest
		.nios2_proc_instruction_master_read             (nios2_proc_instruction_master_read),                          //                                         .read
		.nios2_proc_instruction_master_readdata         (nios2_proc_instruction_master_readdata),                      //                                         .readdata
		.Calibration_s1_address                         (mm_interconnect_0_calibration_s1_address),                    //                           Calibration_s1.address
		.Calibration_s1_write                           (mm_interconnect_0_calibration_s1_write),                      //                                         .write
		.Calibration_s1_readdata                        (mm_interconnect_0_calibration_s1_readdata),                   //                                         .readdata
		.Calibration_s1_writedata                       (mm_interconnect_0_calibration_s1_writedata),                  //                                         .writedata
		.Calibration_s1_chipselect                      (mm_interconnect_0_calibration_s1_chipselect),                 //                                         .chipselect
		.Centaines_s1_address                           (mm_interconnect_0_centaines_s1_address),                      //                             Centaines_s1.address
		.Centaines_s1_readdata                          (mm_interconnect_0_centaines_s1_readdata),                     //                                         .readdata
		.Dizaines_s1_address                            (mm_interconnect_0_dizaines_s1_address),                       //                              Dizaines_s1.address
		.Dizaines_s1_readdata                           (mm_interconnect_0_dizaines_s1_readdata),                      //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.led_s1_address                                 (mm_interconnect_0_led_s1_address),                            //                                   led_s1.address
		.led_s1_write                                   (mm_interconnect_0_led_s1_write),                              //                                         .write
		.led_s1_readdata                                (mm_interconnect_0_led_s1_readdata),                           //                                         .readdata
		.led_s1_writedata                               (mm_interconnect_0_led_s1_writedata),                          //                                         .writedata
		.led_s1_chipselect                              (mm_interconnect_0_led_s1_chipselect),                         //                                         .chipselect
		.Milliers_s1_address                            (mm_interconnect_0_milliers_s1_address),                       //                              Milliers_s1.address
		.Milliers_s1_readdata                           (mm_interconnect_0_milliers_s1_readdata),                      //                                         .readdata
		.nios2_proc_jtag_debug_module_address           (mm_interconnect_0_nios2_proc_jtag_debug_module_address),      //             nios2_proc_jtag_debug_module.address
		.nios2_proc_jtag_debug_module_write             (mm_interconnect_0_nios2_proc_jtag_debug_module_write),        //                                         .write
		.nios2_proc_jtag_debug_module_read              (mm_interconnect_0_nios2_proc_jtag_debug_module_read),         //                                         .read
		.nios2_proc_jtag_debug_module_readdata          (mm_interconnect_0_nios2_proc_jtag_debug_module_readdata),     //                                         .readdata
		.nios2_proc_jtag_debug_module_writedata         (mm_interconnect_0_nios2_proc_jtag_debug_module_writedata),    //                                         .writedata
		.nios2_proc_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_proc_jtag_debug_module_byteenable),   //                                         .byteenable
		.nios2_proc_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_proc_jtag_debug_module_waitrequest),  //                                         .waitrequest
		.nios2_proc_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_proc_jtag_debug_module_debugaccess),  //                                         .debugaccess
		.onchip_memory_s1_address                       (mm_interconnect_0_onchip_memory_s1_address),                  //                         onchip_memory_s1.address
		.onchip_memory_s1_write                         (mm_interconnect_0_onchip_memory_s1_write),                    //                                         .write
		.onchip_memory_s1_readdata                      (mm_interconnect_0_onchip_memory_s1_readdata),                 //                                         .readdata
		.onchip_memory_s1_writedata                     (mm_interconnect_0_onchip_memory_s1_writedata),                //                                         .writedata
		.onchip_memory_s1_byteenable                    (mm_interconnect_0_onchip_memory_s1_byteenable),               //                                         .byteenable
		.onchip_memory_s1_chipselect                    (mm_interconnect_0_onchip_memory_s1_chipselect),               //                                         .chipselect
		.onchip_memory_s1_clken                         (mm_interconnect_0_onchip_memory_s1_clken),                    //                                         .clken
		.Seven_Seg_1_s1_address                         (mm_interconnect_0_seven_seg_1_s1_address),                    //                           Seven_Seg_1_s1.address
		.Seven_Seg_1_s1_write                           (mm_interconnect_0_seven_seg_1_s1_write),                      //                                         .write
		.Seven_Seg_1_s1_readdata                        (mm_interconnect_0_seven_seg_1_s1_readdata),                   //                                         .readdata
		.Seven_Seg_1_s1_writedata                       (mm_interconnect_0_seven_seg_1_s1_writedata),                  //                                         .writedata
		.Seven_Seg_1_s1_chipselect                      (mm_interconnect_0_seven_seg_1_s1_chipselect),                 //                                         .chipselect
		.Seven_Seg_2_s1_address                         (mm_interconnect_0_seven_seg_2_s1_address),                    //                           Seven_Seg_2_s1.address
		.Seven_Seg_2_s1_write                           (mm_interconnect_0_seven_seg_2_s1_write),                      //                                         .write
		.Seven_Seg_2_s1_readdata                        (mm_interconnect_0_seven_seg_2_s1_readdata),                   //                                         .readdata
		.Seven_Seg_2_s1_writedata                       (mm_interconnect_0_seven_seg_2_s1_writedata),                  //                                         .writedata
		.Seven_Seg_2_s1_chipselect                      (mm_interconnect_0_seven_seg_2_s1_chipselect),                 //                                         .chipselect
		.Seven_Seg_3_s1_address                         (mm_interconnect_0_seven_seg_3_s1_address),                    //                           Seven_Seg_3_s1.address
		.Seven_Seg_3_s1_write                           (mm_interconnect_0_seven_seg_3_s1_write),                      //                                         .write
		.Seven_Seg_3_s1_readdata                        (mm_interconnect_0_seven_seg_3_s1_readdata),                   //                                         .readdata
		.Seven_Seg_3_s1_writedata                       (mm_interconnect_0_seven_seg_3_s1_writedata),                  //                                         .writedata
		.Seven_Seg_3_s1_chipselect                      (mm_interconnect_0_seven_seg_3_s1_chipselect),                 //                                         .chipselect
		.Seven_Seg_4_s1_address                         (mm_interconnect_0_seven_seg_4_s1_address),                    //                           Seven_Seg_4_s1.address
		.Seven_Seg_4_s1_write                           (mm_interconnect_0_seven_seg_4_s1_write),                      //                                         .write
		.Seven_Seg_4_s1_readdata                        (mm_interconnect_0_seven_seg_4_s1_readdata),                   //                                         .readdata
		.Seven_Seg_4_s1_writedata                       (mm_interconnect_0_seven_seg_4_s1_writedata),                  //                                         .writedata
		.Seven_Seg_4_s1_chipselect                      (mm_interconnect_0_seven_seg_4_s1_chipselect),                 //                                         .chipselect
		.switcher_s1_address                            (mm_interconnect_0_switcher_s1_address),                       //                              switcher_s1.address
		.switcher_s1_readdata                           (mm_interconnect_0_switcher_s1_readdata),                      //                                         .readdata
		.sysid_1337_control_slave_address               (mm_interconnect_0_sysid_1337_control_slave_address),          //                 sysid_1337_control_slave.address
		.sysid_1337_control_slave_readdata              (mm_interconnect_0_sysid_1337_control_slave_readdata),         //                                         .readdata
		.Unites_s1_address                              (mm_interconnect_0_unites_s1_address),                         //                                Unites_s1.address
		.Unites_s1_readdata                             (mm_interconnect_0_unites_s1_readdata)                         //                                         .readdata
	);

	de1_blinker_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_proc_d_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_proc_jtag_debug_module_reset_reset), // reset_in0.reset
		.clk            (clk_clk),                                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),           // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),       //          .reset_req
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_in1      (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

endmodule
